module sleep (
	input[]
)